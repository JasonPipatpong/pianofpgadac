library verilog;
use verilog.vl_types.all;
entity combine_vlg_vec_tst is
end combine_vlg_vec_tst;
