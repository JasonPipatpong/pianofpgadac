library verilog;
use verilog.vl_types.all;
entity my_I2S_vlg_vec_tst is
end my_I2S_vlg_vec_tst;
